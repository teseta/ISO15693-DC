library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity core_tb is
end core_tb;

architecture sim of core_tb is
    constant CLK_PERIOD : time := 10 ns; -- Periodo del reloj
    
    signal clk_tb : std_logic := '0';
    signal reset_tb : std_logic := '0';
    signal cmd_tb : std_logic := '0';

    component core
        port(
            clk : in std_logic;
            reset : in std_logic;
            cmd : in std_logic
        );
    end component;

begin
    uut: core
    port map (
        clk => clk_tb,
        reset => reset_tb,
        cmd => cmd_tb
    );

    -- Clock generation process
    clk_process: process
    begin
        clk_tb <= '0';
        wait for CLK_PERIOD / 2;
        clk_tb <= '1';
        wait for CLK_PERIOD / 2;
    end process;

    stimulus: process
    begin
        reset_tb <= '1';
        wait for CLK_PERIOD;
        reset_tb <= '0';
        wait for CLK_PERIOD;

        -- Write the first bit then wait for bit period
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
   cmd_tb <= '0';
   wait for 9.44us;
   cmd_tb <= '1';
   wait for 9.44us;
                  
   -- Testing complete
   wait;
    end process;
end sim;

